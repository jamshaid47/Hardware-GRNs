library ieee; 

library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 


entity corr_block is
	port 
		(
		clk			:	in 	std_logic;
		reset	:	in 	std_logic;
		inp1			:	in 	std_logic_vector(15 downto 0);  
		inp2			:	in 	std_logic_vector(15 downto 0);  
		outp1	 :	out 	std_logic_vector (15 downto 0);
		outp2	 :	out 	std_logic_vector (15 downto 0)
		);


	end corr_block ;

architecture behave of corr_block is

type 		data_array18 is array (integer range <>) of std_logic_vector(17 downto 0);

signal  	M 	: 	data_array18(0 to 1023);
signal  	C 	: 	data_array18(0 to 1023);
signal	  sin10, sin20 : std_logic_vector(15 downto 0); 
signal	  sin11, sin21 : std_logic_vector(17 downto 0); 
signal	  sign10, sign20 : std_logic; 
signal   Ms10, Cs10, Cs11 : signed(17 downto 0); 
signal   Ms20, Cs20, Cs21 : signed(17 downto 0); 
signal   outps11, outps21 : signed(35 downto 0); 
signal   outps12, outps22 : signed(23 downto 0); 
signal   addr1, addr2 : unsigned(9 downto 0);  

begin 

--main process that that starts with start of internal clock,
process (reset, clk)
begin
	if (clk'event and clk = '1') then
		if(reset = '0')then
			M <=
			(
			"000000000011011100", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011001", "000000000011011001", "000000000011011001", "000000000011011001",
			"000000000011011001", "000000000011011001", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010110",
			"000000000011010110", "000000000011010110", "000000000011010110", "000000000011010110", "000000000011010110", "000000000011010110", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010100", "000000000011010100",
			"000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011",
			"000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001",
			"000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000",
			"000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111",
			"000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110",
			"000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110",
			"000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110",
			"000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110",
			"000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110",
			"000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001110", "000000000011001111", "000000000011001111",
			"000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111",
			"000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011001111", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000",
			"000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010000", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001", "000000000011010001",
			"000000000011010001", "000000000011010001", "000000000011010001", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010010", "000000000011010011",
			"000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010011", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100",
			"000000000011010100", "000000000011010100", "000000000011010100", "000000000011010100", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010101", "000000000011010110", "000000000011010110",
			"000000000011010110", "000000000011010110", "000000000011010110", "000000000011010110", "000000000011010110", "000000000011010110", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011010111", "000000000011011000",
			"000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011000", "000000000011011001", "000000000011011001", "000000000011011001", "000000000011011001", "000000000011011001", "000000000011011001", "000000000011011001", "000000000011011010", "000000000011011010",
			"000000000011011010", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011010", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011011", "000000000011011100", "000000000011011100", "000000000011011100",
			"000000000011011100", "000000000011011100", "000000000011011100", "000000000011011100", "000000000011011101", "000000000011011101", "000000000011011101", "000000000011011101", "000000000011011101", "000000000011011101", "000000000011011101", "000000000011011110", "000000000011011110", "000000000011011110", "000000000011011110", "000000000011011110",
			"000000000011011110", "000000000011011111", "000000000011011111", "000000000011011111", "000000000011011111", "000000000011011111", "000000000011011111", "000000000011011111", "000000000011100000", "000000000011100000", "000000000011100000", "000000000011100000", "000000000011100000", "000000000011100000", "000000000011100001", "000000000011100001",
			"000000000011100001", "000000000011100001", "000000000011100001", "000000000011100001", "000000000011100010", "000000000011100010", "000000000011100010", "000000000011100010", "000000000011100010", "000000000011100010", "000000000011100011", "000000000011100011", "000000000011100011", "000000000011100011", "000000000011100011", "000000000011100011",
			"000000000011100100", "000000000011100100", "000000000011100100", "000000000011100100", "000000000011100100", "000000000011100100", "000000000011100101", "000000000011100101", "000000000011100101", "000000000011100101", "000000000011100101", "000000000011100101", "000000000011100110", "000000000011100110", "000000000011100110", "000000000011100110",
			"000000000011100110", "000000000011100110", "000000000011100111", "000000000011100111", "000000000011100111", "000000000011100111", "000000000011100111", "000000000011100111", "000000000011101000", "000000000011101000", "000000000011101000", "000000000011101000", "000000000011101000", "000000000011101000", "000000000011101001", "000000000011101001",
			"000000000011101001", "000000000011101001", "000000000011101001", "000000000011101001", "000000000011101010", "000000000011101010", "000000000011101010", "000000000011101010", "000000000011101010", "000000000011101010", "000000000011101010", "000000000011101011", "000000000011101011", "000000000011101011", "000000000011101011", "000000000011101011",
			"000000000011101011", "000000000011101100", "000000000011101100", "000000000011101100", "000000000011101100", "000000000011101100", "000000000011101100", "000000000011101100", "000000000011101101", "000000000011101101", "000000000011101101", "000000000011101101", "000000000011101101", "000000000011101101", "000000000011101101", "000000000011101110",
			"000000000011101110", "000000000011101110", "000000000011101110", "000000000011101110", "000000000011101110", "000000000011101110", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011101111", "000000000011110000",
			"000000000011110000", "000000000011110000", "000000000011110000", "000000000011110000", "000000000011110000", "000000000011110000", "000000000011110000", "000000000011110000", "000000000011110000", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001",
			"000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001",
			"000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001",
			"000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110001", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010",
			"000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110010", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011",
			"000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110011", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110100", "000000000011110101",
			"000000000011110101", "000000000011110101", "000000000011110101", "000000000011110101", "000000000011110101", "000000000011110101", "000000000011110101", "000000000011110101", "000000000011110110", "000000000011110110", "000000000011110110", "000000000011110110", "000000000011110110", "000000000011110110", "000000000011110110", "000000000011110111",
			"000000000011110111", "000000000011110111", "000000000011110111", "000000000011110111", "000000000011110111", "000000000011110111", "000000000011111000", "000000000011111000", "000000000011111000", "000000000011111000", "000000000011111000", "000000000011111000", "000000000011111001", "000000000011111001", "000000000011111001", "000000000011111001",
			"000000000011111001", "000000000011111001", "000000000011111010", "000000000011111010", "000000000011111010", "000000000011111010", "000000000011111010", "000000000011111011", "000000000011111011", "000000000011111011", "000000000011111011", "000000000011111011", "000000000011111100", "000000000011111100", "000000000011111100", "000000000011111100",
			"000000000011111100", "000000000011111101", "000000000011111101", "000000000011111101", "000000000011111101", "000000000011111110", "000000000011111110", "000000000011111110", "000000000011111110", "000000000011111110", "000000000011111111", "000000000011111111", "000000000011111111", "000000000011111111", "000000000100000000", "000000000100000000",
			"000000000100000000", "000000000100000000", "000000000100000001", "000000000100000001", "000000000100000001", "000000000100000001", "000000000100000010", "000000000100000010", "000000000100000010", "000000000100000010", "000000000100000011", "000000000100000011", "000000000100000011", "000000000100000100", "000000000100000100", "000000000100000100",
			"000000000100000100", "000000000100000101", "000000000100000101", "000000000100000101", "000000000100000110", "000000000100000110", "000000000100000110", "000000000100000111", "000000000100000111", "000000000100000111", "000000000100000111", "000000000100001000", "000000000100001000", "000000000100001000", "000000000100001001", "000000000100001001",
			"000000000100001001", "000000000100001010", "000000000100001010", "000000000100001010", "000000000100001011", "000000000100001011", "000000000100001011", "000000000100001100", "000000000100001100", "000000000100001100", "000000000100001101", "000000000100001101", "000000000100001110", "000000000100001110", "000000000100001110", "000000000100001111",
			"000000000100001111", "000000000100001111", "000000000100010000", "000000000100010000", "000000000100010001", "000000000100010001", "000000000100010001", "000000000100010010", "000000000100010010", "000000000100010011", "000000000100010011", "000000000100010011", "000000000100010100", "000000000100010100", "000000000100010101", "000000000100010101",
			"000000000100010110", "000000000100010110", "000000000100010110", "000000000100010111", "000000000100010111", "000000000100011000", "000000000100011000", "000000000100011001", "000000000100011001", "000000000100011010", "000000000100011010", "000000000100011011", "000000000100011011", "000000000100011011", "000000000100011100", "000000000100011100",
			"000000000100011101", "000000000100011101", "000000000100011110", "000000000100011110", "000000000100011111", "000000000100011111", "000000000100100000", "000000000100100000", "000000000100100001", "000000000100100001", "000000000100100010", "000000000100100011", "000000000100100011", "000000000100100100", "000000000100100100", "000000000100100101",
			"000000000100100101", "000000000100100110", "000000000100100110", "000000000100100111", "000000000100101000", "000000000100101000", "000000000100101001", "000000000100101001", "000000000100101010", "000000000100101011", "000000000100101011", "000000000100101100", "000000000100101100", "000000000100101101", "000000000100101110", "000000000100101110",
			"000000000100101111", "000000000100101111", "000000000100110000", "000000000100110001", "000000000100110001", "000000000100110010", "000000000100110011", "000000000100110011", "000000000100110100", "000000000100110101", "000000000100110110", "000000000100110110", "000000000100110111", "000000000100111000", "000000000100111000", "000000000100111001",
			"000000000100111010", "000000000100111010", "000000000100111011", "000000000100111100", "000000000100111101", "000000000100111101", "000000000100111110", "000000000100111111", "000000000101000000", "000000000101000001", "000000000101000001", "000000000101000010", "000000000101000011", "000000000101000100", "000000000101000101", "000000000101000101",
			"000000000101000110", "000000000101000111", "000000000101001000", "000000000101001001", "000000000101001010", "000000000101001011", "000000000101001011", "000000000101001100", "000000000101001101", "000000000101001110", "000000000101001111", "000000000101010000", "000000000101010001", "000000000101010010", "000000000101010011", "000000000101010100",
			"000000000101010101", "000000000101010110", "000000000101010111", "000000000101011000", "000000000101011001", "000000000101011010", "000000000101011011", "000000000101011100", "000000000101011101", "000000000101011110", "000000000101011111", "000000000101100000", "000000000101100001", "000000000101100010", "000000000101100011", "000000000101100100",
			"000000000101100101", "000000000101100111", "000000000101101000", "000000000101101001", "000000000101101010", "000000000101101011", "000000000101101100", "000000000101101110", "000000000101101111", "000000000101110000", "000000000101110001", "000000000101110011", "000000000101110100", "000000000101110101", "000000000101110110", "000000000101111000",
			"000000000101111001", "000000000101111010", "000000000101111100", "000000000101111101", "000000000101111110", "000000000110000000", "000000000110000001", "000000000110000011", "000000000110000100", "000000000110000101", "000000000110000111", "000000000110001000", "000000000110001010", "000000000110001011", "000000000110001101", "000000000110001111",
			"000000000110010000", "000000000110010010", "000000000110010011", "000000000110010101", "000000000110010111", "000000000110011000", "000000000110011010", "000000000110011100", "000000000110011101", "000000000110011111", "000000000110100001", "000000000110100011", "000000000110100100", "000000000110100110", "000000000110101000", "000000000110101010",
			"000000000110101100", "000000000110101110", "000000000110110000", "000000000110110010", "000000000110110100", "000000000110110110", "000000000110111000", "000000000110111010", "000000000110111100", "000000000110111110", "000000000111000000", "000000000111000010", "000000000111000100", "000000000111000111", "000000000111001001", "000000000111001011",
			"000000000111001101", "000000000111010000", "000000000111010010", "000000000111010101", "000000000111010111", "000000000111011010", "000000000111011100", "000000000111011111", "000000000111100001", "000000000111100100", "000000000111100111", "000000000111101001", "000000000111101100", "000000000111101111", "000000000111110010", "000000000111110100",
			"000000000111110111", "000000000111111010", "000000000111111101", "000000001000000000", "000000001000000011", "000000001000000111", "000000001000001010", "000000001000001101", "000000001000010000", "000000001000010100", "000000001000010111", "000000001000011011", "000000001000011110", "000000001000100010", "000000001000100101", "000000001000101001",
			"000000001000101101", "000000001000110001", "000000001000110100", "000000001000111000", "000000001000111100", "000000001001000000", "000000001001000101", "000000001001001001", "000000001001001101", "000000001001010010", "000000001001010110", "000000001001011011", "000000001001011111", "000000001001100100", "000000001001101001", "000000001001101110",
			"000000001001110011", "000000001001111000", "000000001001111101", "000000001010000011", "000000001010001000", "000000001010001110", "000000001010010011", "000000001010011001", "000000001010011111", "000000001010100101", "000000001010101100", "000000001010110010", "000000001010111000", "000000001010111111", "000000001011000110", "000000001011001101",
			"000000001011010100", "000000001011011011", "000000001011100011", "000000001011101010", "000000001011110010", "000000001011111010", "000000001100000011", "000000001100001011", "000000001100010100", "000000001100011101", "000000001100100110", "000000001100101111", "000000001100111001", "000000001101000011", "000000001101001101", "000000001101011000",
			"000000001101100011", "000000001101101110", "000000001101111010", "000000001110000101", "000000001110010010", "000000001110011110", "000000001110101100", "000000001110111001", "000000001111000111", "000000001111010110", "000000001111100101", "000000001111110100", "000000010000000100", "000000010000010101", "000000010000100111", "000000010000111001",
			"000000010001001011", "000000010001011111", "000000010001110011", "000000010010001001", "000000010010011111", "000000010010110110", "000000010011001110", "000000010011100111", "000000010100000010", "000000010100011110", "000000010100111011", "000000010101011010", "000000010101111010", "000000010110011100", "000000010111000001", "000000010111100111",
			"000000011000001111", "000000011000111010", "000000011001101000", "000000011010011001", "000000011011001101", "000000011100000101", "000000011101000001", "000000011110000010", "000000011111001000", "000000100000010100", "000000100001100111", "000000100011000001", "000000100100100100", "000000100110010010", "000000101000001011", "000000101010010010",
			"000000101100101001", "000000101111010101", "000000110010011000", "000000110101111010", "000000111010000000", "000000111110110110", "000001000100101010", "000001001011110010", "000001010100101100", "000001100000001110", "000001110001111100", "000010001000011011", "000010101011000110", "000011101000001010", "000101110011011000", "010010111111111110"
			);
			C <=
			(
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001",
			"000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
			"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111",
			"111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111",
			"111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111111", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110",
			"111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111110", "111111111111111101", "111111111111111101", "111111111111111101",
			"111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101", "111111111111111101",
			"111111111111111101", "111111111111111101", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100",
			"111111111111111100", "111111111111111100", "111111111111111100", "111111111111111100", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011",
			"111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111011", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010",
			"111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111010", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001",
			"111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111001", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000",
			"111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111111000", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111",
			"111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111",
			"111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111",
			"111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111",
			"111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111",
			"111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111", "111111111111110111",
			"111111111111110111", "111111111111110111", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110",
			"111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110110", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101",
			"111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110101", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100", "111111111111110100",
			"111111111111110100", "111111111111110100", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110011", "111111111111110010", "111111111111110010", "111111111111110010", "111111111111110010", "111111111111110010",
			"111111111111110010", "111111111111110010", "111111111111110010", "111111111111110010", "111111111111110001", "111111111111110001", "111111111111110001", "111111111111110001", "111111111111110001", "111111111111110001", "111111111111110001", "111111111111110001", "111111111111110000", "111111111111110000", "111111111111110000", "111111111111110000",
			"111111111111110000", "111111111111110000", "111111111111110000", "111111111111101111", "111111111111101111", "111111111111101111", "111111111111101111", "111111111111101111", "111111111111101111", "111111111111101111", "111111111111101110", "111111111111101110", "111111111111101110", "111111111111101110", "111111111111101110", "111111111111101110",
			"111111111111101101", "111111111111101101", "111111111111101101", "111111111111101101", "111111111111101101", "111111111111101101", "111111111111101100", "111111111111101100", "111111111111101100", "111111111111101100", "111111111111101100", "111111111111101011", "111111111111101011", "111111111111101011", "111111111111101011", "111111111111101011",
			"111111111111101010", "111111111111101010", "111111111111101010", "111111111111101010", "111111111111101010", "111111111111101001", "111111111111101001", "111111111111101001", "111111111111101001", "111111111111101001", "111111111111101000", "111111111111101000", "111111111111101000", "111111111111101000", "111111111111100111", "111111111111100111",
			"111111111111100111", "111111111111100111", "111111111111100110", "111111111111100110", "111111111111100110", "111111111111100110", "111111111111100101", "111111111111100101", "111111111111100101", "111111111111100101", "111111111111100100", "111111111111100100", "111111111111100100", "111111111111100100", "111111111111100011", "111111111111100011",
			"111111111111100011", "111111111111100010", "111111111111100010", "111111111111100010", "111111111111100010", "111111111111100001", "111111111111100001", "111111111111100001", "111111111111100000", "111111111111100000", "111111111111100000", "111111111111100000", "111111111111011111", "111111111111011111", "111111111111011111", "111111111111011110",
			"111111111111011110", "111111111111011110", "111111111111011101", "111111111111011101", "111111111111011101", "111111111111011100", "111111111111011100", "111111111111011100", "111111111111011011", "111111111111011011", "111111111111011010", "111111111111011010", "111111111111011010", "111111111111011001", "111111111111011001", "111111111111011001",
			"111111111111011000", "111111111111011000", "111111111111010111", "111111111111010111", "111111111111010111", "111111111111010110", "111111111111010110", "111111111111010101", "111111111111010101", "111111111111010101", "111111111111010100", "111111111111010100", "111111111111010011", "111111111111010011", "111111111111010010", "111111111111010010",
			"111111111111010010", "111111111111010001", "111111111111010001", "111111111111010000", "111111111111010000", "111111111111001111", "111111111111001111", "111111111111001110", "111111111111001110", "111111111111001101", "111111111111001101", "111111111111001100", "111111111111001100", "111111111111001011", "111111111111001011", "111111111111001010",
			"111111111111001010", "111111111111001001", "111111111111001001", "111111111111001000", "111111111111001000", "111111111111000111", "111111111111000110", "111111111111000110", "111111111111000101", "111111111111000101", "111111111111000100", "111111111111000100", "111111111111000011", "111111111111000010", "111111111111000010", "111111111111000001",
			"111111111111000001", "111111111111000000", "111111111110111111", "111111111110111111", "111111111110111110", "111111111110111101", "111111111110111101", "111111111110111100", "111111111110111011", "111111111110111011", "111111111110111010", "111111111110111001", "111111111110111001", "111111111110111000", "111111111110110111", "111111111110110110",
			"111111111110110110", "111111111110110101", "111111111110110100", "111111111110110011", "111111111110110011", "111111111110110010", "111111111110110001", "111111111110110000", "111111111110110000", "111111111110101111", "111111111110101110", "111111111110101101", "111111111110101100", "111111111110101011", "111111111110101011", "111111111110101010",
			"111111111110101001", "111111111110101000", "111111111110100111", "111111111110100110", "111111111110100101", "111111111110100100", "111111111110100011", "111111111110100010", "111111111110100001", "111111111110100000", "111111111110011111", "111111111110011110", "111111111110011101", "111111111110011100", "111111111110011011", "111111111110011010",
			"111111111110011001", "111111111110011000", "111111111110010111", "111111111110010110", "111111111110010101", "111111111110010100", "111111111110010011", "111111111110010010", "111111111110010000", "111111111110001111", "111111111110001110", "111111111110001101", "111111111110001100", "111111111110001010", "111111111110001001", "111111111110001000",
			"111111111110000111", "111111111110000101", "111111111110000100", "111111111110000011", "111111111110000001", "111111111110000000", "111111111101111111", "111111111101111101", "111111111101111100", "111111111101111010", "111111111101111001", "111111111101111000", "111111111101110110", "111111111101110101", "111111111101110011", "111111111101110001",
			"111111111101110000", "111111111101101110", "111111111101101101", "111111111101101011", "111111111101101001", "111111111101101000", "111111111101100110", "111111111101100100", "111111111101100010", "111111111101100001", "111111111101011111", "111111111101011101", "111111111101011011", "111111111101011001", "111111111101010111", "111111111101010101",
			"111111111101010100", "111111111101010010", "111111111101001111", "111111111101001101", "111111111101001011", "111111111101001001", "111111111101000111", "111111111101000101", "111111111101000011", "111111111101000000", "111111111100111110", "111111111100111100", "111111111100111001", "111111111100110111", "111111111100110101", "111111111100110010",
			"111111111100110000", "111111111100101101", "111111111100101010", "111111111100101000", "111111111100100101", "111111111100100010", "111111111100011111", "111111111100011101", "111111111100011010", "111111111100010111", "111111111100010100", "111111111100010001", "111111111100001110", "111111111100001011", "111111111100000111", "111111111100000100",
			"111111111100000001", "111111111011111101", "111111111011111010", "111111111011110110", "111111111011110011", "111111111011101111", "111111111011101100", "111111111011101000", "111111111011100100", "111111111011100000", "111111111011011100", "111111111011011000", "111111111011010100", "111111111011001111", "111111111011001011", "111111111011000111",
			"111111111011000010", "111111111010111101", "111111111010111001", "111111111010110100", "111111111010101111", "111111111010101010", "111111111010100101", "111111111010011111", "111111111010011010", "111111111010010100", "111111111010001111", "111111111010001001", "111111111010000011", "111111111001111101", "111111111001110111", "111111111001110000",
			"111111111001101010", "111111111001100011", "111111111001011100", "111111111001010101", "111111111001001110", "111111111001000110", "111111111000111111", "111111111000110111", "111111111000101111", "111111111000100110", "111111111000011110", "111111111000010101", "111111111000001100", "111111111000000011", "111111110111111001", "111111110111101111",
			"111111110111100101", "111111110111011011", "111111110111010000", "111111110111000101", "111111110110111001", "111111110110101101", "111111110110100001", "111111110110010100", "111111110110000111", "111111110101111001", "111111110101101011", "111111110101011100", "111111110101001101", "111111110100111101", "111111110100101100", "111111110100011011",
			"111111110100001001", "111111110011110111", "111111110011100011", "111111110011001111", "111111110010111010", "111111110010100100", "111111110010001101", "111111110001110100", "111111110001011011", "111111110001000000", "111111110000100100", "111111110000000110", "111111101111100111", "111111101111000110", "111111101110100011", "111111101101111110",
			"111111101101010111", "111111101100101101", "111111101100000001", "111111101011010001", "111111101010011110", "111111101001101000", "111111101000101101", "111111100111101110", "111111100110101010", "111111100101100000", "111111100100001111", "111111100010110110", "111111100001010101", "111111011111101010", "111111011101110011", "111111011011101110",
			"111111011001011001", "111111010110110000", "111111010011101111", "111111010000010001", "111111001100001101", "111111000111011011", "111111000001101010", "111110111010100111", "111110110001110001", "111110100110010101", "111110010100110100", "111101111110011100", "111101011011111010", "111100011111000010", "111010010100000101", "101101001000001010"
			);


			else
			--Cycle 0
			if(inp1(15) = '0')then
				addr1 <= unsigned(inp1(14 downto 5));
				sign10 <= '0';
  			else
				addr1 <= unsigned(not(inp1(14 downto 5)));
				sign10 <= '1';
			end if;
			sin10 <= inp1;
			
			if(inp2(15) = '0')then
				addr2 <= unsigned(inp2(14 downto 5));
				sign20 <= '0';
  			else
				addr2 <= unsigned(not(inp2(14 downto 5)));
				sign20 <= '1';
			end if;
			sin20 <= inp2;
			
			--Cycle 1
			if(sign10 = '0')then
				Ms10 <= signed(M(to_integer(addr1)));
				Cs10 <= signed(C(to_integer(addr1)));
  			else
				Ms10 <= signed(M(to_integer(addr1)));
				Cs10 <= -signed(C(to_integer(addr1)));
			end if;
			sin11 <= sin10(15) & sin10(15) & sin10;--5.13
			
			if(sign20 = '0')then
				Ms20 <= signed(M(to_integer(addr2)));
				Cs20 <= signed(C(to_integer(addr2)));
  			else
				Ms20 <= signed(M(to_integer(addr2)));
				Cs20 <= -signed(C(to_integer(addr2)));
			end if;
			sin21 <= sin20(15) & sin20(15) & sin20;--5.13
			
			--Cycle 2
			outps11 <= Ms10*signed(sin11);--10.8*5.13=15.21
			Cs11 <= Cs10; --12.6

			outps21 <= Ms20*signed(sin21);--10.8*5.13=15.21
			Cs21 <= Cs20; --12.6

			--Cycle 3
			outps12 <= (outps11(32 downto 9)) + (Cs11 & "000000"); --12.12 + 12.12
			outps22 <= (outps21(32 downto 9)) + (Cs21 & "000000"); --12.12 + 12.12
		end if;
	end if;
end process ;
			outp1 <= std_logic_vector(outps12(15 downto 0));
			outp2 <= std_logic_vector(outps22(15 downto 0));
end behave;








		

